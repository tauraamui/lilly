module ui
