module draw

fn new_context() Contextable {
	return Context{}
}

