// Copyright 2025 The Lilly Edtior contributors
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

module clipboardv3

fn test_linux_clipboard_sets_contents() {
	mut lc := new_linux_clipboard()
	defer { lc.set_content(ClipboardContent{}) }

	lc.set_content(ClipboardContent{ data: "this is a test line of text" })
	assert lc.get_content()! == ClipboardContent{
		data: "this is a test line of text"
	}
}

fn test_linux_clipboard_via_interface_sets_contents() {
	mut c := new()
	defer { c.set_content(ClipboardContent{}) }

	c.set_content(ClipboardContent{ data: "this is a test line of text via interface wrap" })
	assert c.get_content()! == ClipboardContent{
		data: "this is a test line of text via interface wrap"
	}
}

