// Copyright 2024 The Lilly Editor contributors
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

module clipboardv2

pub enum ContentType as u8 {
	@none
	inline
	block
}

pub struct ClipboardContent {
pub:
	type        ContentType
	data         string
}

pub struct Clipboard {
mut:
	content ClipboardContent
}

pub fn new() &Clipboard {
	return &Clipboard{
		content: ClipboardContent{ type: .none }
	}
}

pub fn (mut clipboard Clipboard) get_content() ClipboardContent {
	return clipboard.content
}

pub fn (mut clipboard Clipboard) set_content(content ClipboardContent) {
	clipboard.content = content
	// update system clipboard here
}
