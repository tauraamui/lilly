module ui

struct TodoCommentPickerModal {
}
