// Copyright 2024 The Lilly Editor contributors
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

module clipboard

@[heap]
struct MockClipboard {
mut:
	copied_content        string
	was_copy_unsuccessful bool
}

fn (mut mockclipboard MockClipboard) copy(text string) bool {
	mockclipboard.copied_content = text
	return !mockclipboard.was_copy_unsuccessful
}

fn (mut mockclipboard MockClipboard) paste() string {
	return mockclipboard.copied_content
}
