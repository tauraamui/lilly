module main

import lib.utf8

fn main() {
	println(utf8.emojis)
}

