module main

pub const emoji_shark_char = "🦈"

