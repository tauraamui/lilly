module ui

pub struct BufferEditor {}
