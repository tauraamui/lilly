module main

fn main() {
	println(emojis)
}

