module draw

import term.ui as tui

struct Grid {
	data []Cell
}

fn (mut grid Grid) set_cell(x int, y int, c Cell) {
}

struct Cell {
	data     ?rune
	fg_color Color
	bg_color Color
}

struct ImmediateContext {
	render_debug bool
mut:
	ref            &tui.Context
	previous_frame Grid
	frame          Grid
}

type Runner = fn () !

pub fn new_immediate_context(cfg Config) (&Contextable, Runner) {
	ctx := ImmediateContext{
		render_debug: cfg.render_debug
		ref: tui.init(
			user_data: cfg.user_data
			event_fn:  fn [cfg] (e &tui.Event, app voidptr) {
				cfg.event_fn(Event{e}, app)
			}
			frame_fn:             cfg.frame_fn
			capture_events:       cfg.capture_events
			use_alternate_buffer: cfg.use_alternate_buffer
			frame_rate: 30
		)
	}
	return ctx, unsafe { ctx.run }
}

fn (mut ctx ImmediateContext) rate_limit_draws() bool {
	return true
}

fn (mut ctx ImmediateContext) render_debug() bool { return ctx.render_debug }

fn (mut ctx ImmediateContext) window_width() int {
	return 100
}

fn (mut ctx ImmediateContext) window_height() int {
	return 100
}

fn (mut ctx ImmediateContext) set_cursor_position(x int, y int) {
	ctx.ref.set_cursor_position(x, y)
}

fn (mut ctx ImmediateContext) show_cursor() {
	ctx.ref.show_cursor()
}

fn (mut ctx ImmediateContext) hide_cursor() {
	ctx.ref.hide_cursor()
}

fn (mut ctx ImmediateContext) draw_text(x int, y int, text string) {
	for c_char in text.runes() {
	}
	ctx.ref.draw_text(x, y, text)
}

fn (mut ctx ImmediateContext) write(c string) {
	ctx.ref.write(c)
}

fn (mut ctx ImmediateContext) draw_rect(x int, y int, width int, height int) {
	ctx.ref.draw_rect(x, y, x + (width - 1), y + (height - 1))
}

fn (mut ctx ImmediateContext) draw_point(x int, y int) {
	ctx.ref.draw_point(x, y)
}

fn (mut ctx ImmediateContext) bold() {
	ctx.ref.bold()
}

fn (mut ctx ImmediateContext) set_color(c Color) {
	ctx.ref.set_color(tui.Color{ r: c.r, g: c.g, b: c.b })
}

fn (mut ctx ImmediateContext) set_bg_color(c Color) {
	ctx.ref.set_bg_color(tui.Color{ r: c.r, g: c.g, b: c.b })
}

fn (mut ctx ImmediateContext) reset_color() {
	ctx.ref.reset_color()
}

fn (mut ctx ImmediateContext) reset_bg_color() {
	ctx.ref.reset_bg_color()
}

fn (mut ctx ImmediateContext) reset() {
	ctx.ref.reset()
}

fn (mut ctx ImmediateContext) run() ! {
	return ctx.ref.run()
}

fn (mut ctx ImmediateContext) clear() {
	ctx.ref.clear()
}

fn (mut ctx ImmediateContext) flush() {
	ctx.ref.flush()
}

