module workspace

pub struct Workspace {
}

pub fn open_workspace(root_path string) !Workspace {
	return error("workspace not implemented yet")
}

