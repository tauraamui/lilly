module draw

fn test_new_immediate_mode_ctx() {
	ctx, run := new_immediate_context(
		render_debug: false
	)
}


