module utf8

const emoji_shark_char = "🦈"
