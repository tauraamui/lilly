module clipboard
