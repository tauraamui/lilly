module utf8

pub const emoji_shark_char = "🦈"

pub const emojis = {
	"shark": "🦈"
	"whale": "🐳"
	"dolphin": "🐬"
	"octopus": "🐙"
	"crab": "🦀"
	"squid": "🦑"
	"turtle": "🐢"
	"fish": "🐟"
	"tropical_fish": "🐠"
	"blowfish": "🐡"
	"seal": "🦭"
	"diving_mask": "🤿"
}
