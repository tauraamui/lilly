module main

fn main() {
	println(emoji_shark_char)
}

