module utf8

pub const emoji_shark_char = '🦈'
