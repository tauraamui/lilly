// Copyright 2025 The Lilly Editor contributors
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

module draw

@[params]
pub struct PaintShapeTextArgs {
pub:
	x        int
	y        int
	fg_color Color
	text     string
}

pub fn paint_shape_text(mut ctx Contextable, x int, y int, color Color, text string) {
	ctx.set_color(r: color.r, g: color.g, b: color.b)
	ctx.reset_bg_color()
	ctx.draw_text(x, y, text)
}

@[params]
pub struct PaintTextOnBackgroundArgs {
pub:
	x int
	y int
	bg_color Color
	fg_color Color
	text     string
}

pub fn paint_text_on_background(mut ctx Contextable, args PaintTextOnBackgroundArgs) {
// pub fn paint_text_on_background(mut ctx Contextable, x int, y int, bg_color Color, fg_color Color, text string) {
	bg_color := args.bg_color
	fg_color := args.fg_color
	ctx.set_bg_color(r: bg_color.r, g: bg_color.g, b: bg_color.b)
	ctx.set_color(r: fg_color.r, g: fg_color.g, b: fg_color.b)
	ctx.draw_text(args.x, args.y, args.text)
}
