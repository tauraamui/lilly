module clipboardv3

fn test_clipboard_native_implementation() {
	ct := ContentType.inline
}

