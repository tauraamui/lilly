// Copyright 2025 The Lilly Editor contributors
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

module clipboard

import clipboard as stdlib_clipboard
import os

fn new_clipboard() Clipboard {
	// NOTE(tauraamui): temp disable wayland clipboard support
	// if os_running_wayland() {
	// 	$if !test { return WaylandClipboard{} }
	// }
	$if test {
		return MockClipboard{}
	}
	return StdLibClipboard{
		ref: stdlib_clipboard.new_primary()
	}
}

fn os_running_wayland() bool {
	return os.getenv('WAYLAND_DISPLAY').len > 0
}
