module workspace

pub struct Syntax {
pub:
	name       string
	extensions []string
	keywords   []string
	literals   []string
}

